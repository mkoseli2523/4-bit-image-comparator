f4
.lib '/class/ece482/gpdk045_mos' TT
.param TCK = 0.4n
.param trf_ck = 5p
.param CK_pw = 0.5*TCK

** Library name: final_v2
** Cell name: register_2
** View name: schematic
.subckt register_2 clk clk_bar d q rst vdd vss
mpm3 net4 x vdd vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm2 q clk_bar net4 vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm1 x clk net2 vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm0 net2 d vdd vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mnm17 q rst vss vss g45n1svt L=45e-9 W=5.76e-6 AD='5.76e-6/ceil(575.9995e-3)<119.5e-9?(floor(ceil(575.9995e-3)/2.0)*(14.4e-15+(5.76e-6/ceil(575.9995e-3))*100e-9)+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9:0))/1:(floor(ceil(575.9995e-3)/2.0)*(110e-9*(5.76e-6/ceil(575.9995e-3)))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?140e-9*(5.76e-6/ceil(575.9995e-3)):0))/1' AS='5.76e-6/ceil(575.9995e-3)<119.5e-9?(((14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9)+floor((ceil(575.9995e-3)-1)/2.0)*(14.4e-15+(5.76e-6/ceil(575.9995e-3))*100e-9))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9:0))/1:((140e-9*(5.76e-6/ceil(575.9995e-3))+floor((ceil(575.9995e-3)-1)/2.0)*(110e-9*(5.76e-6/ceil(575.9995e-3))))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?140e-9*(5.76e-6/ceil(575.9995e-3)):0))/1'
+PD='5.76e-6/ceil(575.9995e-3)<119.5e-9?(floor(ceil(575.9995e-3)/2.0)*680e-9+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(575.9995e-3)/2.0)*(220e-9+2*(5.76e-6/ceil(575.9995e-3)))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?280e-9+2*(5.76e-6/ceil(575.9995e-3)):0))/1' PS='5.76e-6/ceil(575.9995e-3)<119.5e-9?((580e-9+floor((ceil(575.9995e-3)-1)/2.0)*680e-9)+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(5.76e-6/ceil(575.9995e-3)))+floor((ceil(575.9995e-3)-1)/2.0)*(220e-9+2*(5.76e-6/ceil(575.9995e-3))))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?280e-9+2*(5.76e-6/ceil(575.9995e-3)):0))/1'
+NRD='5.76e-6/ceil(575.9995e-3)<119.5e-9?(floor(ceil(575.9995e-3)/2.0)*(14.4e-15+(5.76e-6/ceil(575.9995e-3))*100e-9)+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9:0))/1:((floor(ceil(575.9995e-3)/2.0)*(110e-9*(5.76e-6/ceil(575.9995e-3)))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)!=0?140e-9*(5.76e-6/ceil(575.9995e-3)):0))/1)/((((5.76e-6/ceil(575.9995e-3))*ceil(575.9995e-3))*(5.76e-6/ceil(575.9995e-3)))*ceil(575.9995e-3))'
+NRS='5.76e-6/ceil(575.9995e-3)<119.5e-9?(((14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9)+floor((ceil(575.9995e-3)-1)/2.0)*(14.4e-15+(5.76e-6/ceil(575.9995e-3))*100e-9))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?14.4e-15+(5.76e-6/ceil(575.9995e-3))*50e-9:0))/1:(((140e-9*(5.76e-6/ceil(575.9995e-3))+floor((ceil(575.9995e-3)-1)/2.0)*(110e-9*(5.76e-6/ceil(575.9995e-3))))+(ceil(575.9995e-3)/2-floor(ceil(575.9995e-3)/2)==0?140e-9*(5.76e-6/ceil(575.9995e-3)):0))/1)/((((5.76e-6/ceil(575.9995e-3))*ceil(575.9995e-3))*(5.76e-6/ceil(575.9995e-3)))*ceil(575.9995e-3))' M=1
mnm3 net3 x vss vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm2 q clk net3 vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm1 net1 d vss vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm0 x clk_bar net1 vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
c5 clk vss 2e-15
c4 clk_bar vss 2e-15
c3 clk vss 2e-15
c2 clk_bar vss 2e-15
c1 x vss 2e-15
c0 d vss 2e-15
c11 rst vss 2e-15
.ends register_2
** End of subcircuit definition.

** Library name: final_v2
** Cell name: inv
** View name: schematic
.subckt inv vdd vss in out
mpm0 out in vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm0 out in vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends inv
** End of subcircuit definition.

** Library name: final_v2
** Cell name: clk_deskew
** View name: schematic
.subckt clk_deskew ck ck_bar clk vdd vss
mnm5 ck clk_out vss vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm4 clk_out clk vss vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm1 ck_bar t_out vss vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mnm0 t_out vdd clk vss g45n1svt L=45e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mpm5 ck clk_out vdd vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm4 clk_out clk vdd vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm1 ck_bar t_out vdd vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
mpm0 t_out vss clk vdd g45p1svt L=45e-9 W=960e-9 AD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1' AS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1'
+PD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*680e-9+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(95.9995e-3)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1' PS='960e-9/ceil(95.9995e-3)<119.5e-9?((580e-9+floor((ceil(95.9995e-3)-1)/2.0)*680e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(960e-9/ceil(95.9995e-3)))+floor((ceil(95.9995e-3)-1)/2.0)*(220e-9+2*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?280e-9+2*(960e-9/ceil(95.9995e-3)):0))/1'
+NRD='960e-9/ceil(95.9995e-3)<119.5e-9?(floor(ceil(95.9995e-3)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9)+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:((floor(ceil(95.9995e-3)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3)))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)!=0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' NRS='960e-9/ceil(95.9995e-3)<119.5e-9?(((14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9)+floor((ceil(95.9995e-3)-1)/2.0)*(14.4e-15+(960e-9/ceil(95.9995e-3))*100e-9))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?14.4e-15+(960e-9/ceil(95.9995e-3))*50e-9:0))/1:(((140e-9*(960e-9/ceil(95.9995e-3))+floor((ceil(95.9995e-3)-1)/2.0)*(110e-9*(960e-9/ceil(95.9995e-3))))+(ceil(95.9995e-3)/2-floor(ceil(95.9995e-3)/2)==0?140e-9*(960e-9/ceil(95.9995e-3)):0))/1)/((((960e-9/ceil(95.9995e-3))*ceil(95.9995e-3))*(960e-9/ceil(95.9995e-3)))*ceil(95.9995e-3))' M=1
.ends clk_deskew
** End of subcircuit definition.

** Library name: final_v2
** Cell name: f4v2
** View name: schematic
xi1 net4 net1 net5 q rst vdd vss register_2
xi0 net6 net2 net1 net4 rst vdd vss register_2
xi3 vdd vss q net5 inv
xi2 vdd vss net4 net1 inv
xi4 net6 net2 clk vdd vss clk_deskew

vclk clk 0 pulse(0 1.1 trf_ck trf_ck trf_ck CK_pw TCK)

vVDD vdd 0 1.1
vVSS vss 0 0

.tran 0.1ps 20ns

.option post
.end
